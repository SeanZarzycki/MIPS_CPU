library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity id_ex_reg is

end id_ex_reg;

architecture beh of id_ex_reg is

begin

end beh;