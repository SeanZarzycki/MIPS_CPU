library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity if_id_reg is

end if_id_reg;

architecture beh of if_id_reg is

begin

end beh;